module ALU_4_Bit(input a,input b,output reg )


endmodule