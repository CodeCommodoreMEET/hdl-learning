module endmodule 